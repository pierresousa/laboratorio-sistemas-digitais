library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity tb_centro_recebimento_graos is

end tb_centro_recebimento_graos;


architecture teste of tb_centro_recebimento_graos is

component centro_recebimento_graos is 
port (
        RESET   : in    std_logic; -- reset input
        CLOCK   : in    std_logic; -- clock input
		PODE_PESAR       : in    std_logic; -- permite pesagem do caminhao
		PESO_BRUTO       : in    std_logic_vector(28 downto 0); -- peso bruto do caminhao com carga
		PESO_CAMINHAO       : in    std_logic_vector(28 downto 0); -- peso bruto do caminhao somente
		TIPO_GRAO       : in    std_logic_vector(1 downto 0); -- informa o tipo do grao
		LOCAL_SILO       : out    std_logic_vector(1 downto 0); -- informa o silo referente ao grao
		SENSOR_VAGA_SOJA       : in    std_logic; -- verifica se o silo de soja esta ocupado
		LAMPADA_VAGA_SOJA       : out    std_logic; -- informa se o silo de soja esta ocupado
		SENSOR_VAGA_ARROZ       : in    std_logic; -- verifica se o silo de arroz esta ocupado
		LAMPADA_VAGA_ARROZ       : out    std_logic; -- informa se o silo de arroz esta ocupado
		SENSOR_VAGA_FEIJAO       : in    std_logic; -- verifica se o silo de feijao esta ocupado
		LAMPADA_VAGA_FEIJAO       : out    std_logic; -- informa se o silo de feijao esta ocupado
		MOTOR_ESCOTILHA_SOJA       : out    std_logic_vector(1 downto 0); -- abre a escotilha do silo soja
		MOTOR_ESCOTILHA_ARROZ       : out    std_logic_vector(1 downto 0); -- abre a escotilha do silo arroz
		MOTOR_ESCOTILHA_FEIJAO       : out    std_logic_vector(1 downto 0); -- abre a escotilha do silo feijao
		PESO_CARGA       : out    std_logic_vector(28 downto 0); -- peso da carga
		VALOR_CARGA       : out    std_logic_vector(31 downto 0) -- valor a ser pago pela carga
);
end component;

signal CLOCK, RESET, PODE_PESAR, SENSOR_VAGA_SOJA, LAMPADA_VAGA_SOJA, SENSOR_VAGA_ARROZ, LAMPADA_VAGA_ARROZ, SENSOR_VAGA_FEIJAO, LAMPADA_VAGA_FEIJAO: std_logic;
signal PESO_BRUTO, PESO_CAMINHAO, PESO_CARGA: std_logic_vector(28 downto 0);
signal VALOR_CARGA: std_logic_vector(31 downto 0);
signal TIPO_GRAO, LOCAL_SILO, MOTOR_ESCOTILHA_SOJA, MOTOR_ESCOTILHA_ARROZ, MOTOR_ESCOTILHA_FEIJAO: std_logic_vector(1 downto 0);
begin
instancia_centro_recebimento_graos: centro_recebimento_graos port map (CLOCK=>CLOCK,
																							  RESET=>RESET,
																							  PODE_PESAR=>PODE_PESAR,
																							  PESO_BRUTO=>PESO_BRUTO,
																							  PESO_CAMINHAO=>PESO_CAMINHAO,
																							  TIPO_GRAO=>TIPO_GRAO,
																							  LOCAL_SILO=>LOCAL_SILO,
																							  SENSOR_VAGA_SOJA=>SENSOR_VAGA_SOJA,
																							  SENSOR_VAGA_ARROZ=>SENSOR_VAGA_ARROZ,
																							  SENSOR_VAGA_FEIJAO=>SENSOR_VAGA_FEIJAO,
																							  LAMPADA_VAGA_SOJA=>LAMPADA_VAGA_SOJA,
																							  LAMPADA_VAGA_ARROZ=>LAMPADA_VAGA_ARROZ,
																							  LAMPADA_VAGA_FEIJAO=>LAMPADA_VAGA_FEIJAO,
																							  MOTOR_ESCOTILHA_SOJA=>MOTOR_ESCOTILHA_SOJA,
																							  MOTOR_ESCOTILHA_ARROZ=>MOTOR_ESCOTILHA_ARROZ,
																							  MOTOR_ESCOTILHA_FEIJAO=>MOTOR_ESCOTILHA_FEIJAO,
																							  PESO_CARGA=>PESO_CARGA,
																							  VALOR_CARGA=>VALOR_CARGA);
CLOCK <= '0',
			'1' after 5 ns, '0' after 10 ns, 
			'1' after 15 ns, '0' after 20 ns, 
			'1' after 25 ns, '0' after 30 ns, 
			'1' after 35 ns, '0' after 40 ns, 
			'1' after 45 ns, '0' after 50 ns, 
			'1' after 55 ns, '0' after 60 ns, 
			'1' after 65 ns, '0' after 70 ns, 
			'1' after 75 ns, '0' after 80 ns,
			'1' after 85 ns, '0' after 90 ns,
			'1' after 95 ns, '0' after 100 ns,
			'1' after 105 ns, '0' after 110 ns, 
			'1' after 115 ns, '0' after 120 ns, 
			'1' after 125 ns, '0' after 130 ns, 
			'1' after 135 ns, '0' after 140 ns, 
			'1' after 145 ns, '0' after 150 ns, 
			'1' after 155 ns, '0' after 160 ns, 
			'1' after 165 ns, '0' after 170 ns, 
			'1' after 175 ns, '0' after 180 ns,
			'1' after 185 ns, '0' after 190 ns,
			'1' after 195 ns, '0' after 200 ns,
			'1' after 205 ns, '0' after 210 ns, 
			'1' after 215 ns, '0' after 220 ns, 
			'1' after 225 ns, '0' after 230 ns, 
			'1' after 235 ns, '0' after 240 ns, 
			'1' after 245 ns, '0' after 250 ns, 
			'1' after 255 ns, '0' after 260 ns, 
			'1' after 265 ns, '0' after 270 ns, 
			'1' after 275 ns, '0' after 280 ns,
			'1' after 285 ns, '0' after 290 ns,
			'1' after 295 ns, '0' after 300 ns,
			'1' after 305 ns, '0' after 310 ns, 
			'1' after 315 ns, '0' after 320 ns, 
			'1' after 325 ns, '0' after 330 ns, 
			'1' after 335 ns, '0' after 340 ns, 
			'1' after 345 ns, '0' after 350 ns, 
			'1' after 355 ns, '0' after 360 ns, 
			'1' after 365 ns, '0' after 370 ns, 
			'1' after 375 ns, '0' after 380 ns,
			'1' after 385 ns, '0' after 390 ns,
			'1' after 395 ns, '0' after 400 ns,
			'1' after 405 ns, '0' after 410 ns, 
			'1' after 415 ns, '0' after 420 ns, 
			'1' after 425 ns, '0' after 430 ns, 
			'1' after 435 ns, '0' after 440 ns, 
			'1' after 445 ns, '0' after 450 ns, 
			'1' after 455 ns, '0' after 460 ns, 
			'1' after 465 ns, '0' after 470 ns, 
			'1' after 475 ns, '0' after 480 ns,
			'1' after 485 ns, '0' after 490 ns,
			'1' after 495 ns, '0' after 500 ns,
			'1' after 505 ns, '0' after 510 ns, 
			'1' after 515 ns, '0' after 520 ns, 
			'1' after 525 ns, '0' after 530 ns, 
			'1' after 535 ns, '0' after 540 ns, 
			'1' after 545 ns, '0' after 550 ns, 
			'1' after 555 ns, '0' after 560 ns, 
			'1' after 565 ns, '0' after 570 ns, 
			'1' after 575 ns, '0' after 580 ns,
			'1' after 585 ns, '0' after 590 ns,
			'1' after 595 ns, '0' after 600 ns,
			'1' after 605 ns, '0' after 610 ns, 
			'1' after 615 ns, '0' after 620 ns, 
			'1' after 625 ns, '0' after 630 ns, 
			'1' after 635 ns, '0' after 640 ns, 
			'1' after 645 ns, '0' after 650 ns, 
			'1' after 655 ns, '0' after 660 ns, 
			'1' after 665 ns, '0' after 670 ns, 
			'1' after 675 ns, '0' after 680 ns,
			'1' after 685 ns, '0' after 690 ns,
			'1' after 695 ns, '0' after 700 ns,
			'1' after 705 ns, '0' after 710 ns, 
			'1' after 715 ns, '0' after 720 ns, 
			'1' after 725 ns, '0' after 730 ns, 
			'1' after 735 ns, '0' after 740 ns, 
			'1' after 745 ns, '0' after 750 ns, 
			'1' after 755 ns, '0' after 760 ns, 
			'1' after 765 ns, '0' after 770 ns, 
			'1' after 775 ns, '0' after 780 ns,
			'1' after 785 ns, '0' after 790 ns,
			'1' after 795 ns, '0' after 800 ns;
RESET <= '1',
			'0' after 4 ns;
PODE_PESAR <= '0', 
		'1' after 4 ns, '0' after 10 ns, 
		'1' after 24 ns, '0' after 30 ns, 
		'1' after 44 ns, '0' after 50 ns, 
		'1' after 64 ns, '0' after 70 ns, 
		'1' after 84 ns, '0' after 90 ns,
		'1' after 104 ns, '0' after 110 ns, 
		'1' after 124 ns, '0' after 130 ns,  
		'1' after 144 ns, '0' after 150 ns, 
		'1' after 164 ns, '0' after 170 ns, 
		'1' after 184 ns, '0' after 190 ns,
		'1' after 204 ns, '0' after 210 ns,  
		'1' after 224 ns, '0' after 230 ns, 
		'1' after 244 ns, '0' after 250 ns, 
		'1' after 264 ns, '0' after 270 ns, 
		'1' after 284 ns, '0' after 290 ns,
		'1' after 304 ns, '0' after 310 ns,  
		'1' after 324 ns, '0' after 330 ns, 
		'1' after 344 ns, '0' after 350 ns,  
		'1' after 364 ns, '0' after 370 ns, 
		'1' after 384 ns, '0' after 390 ns,
		'1' after 404 ns, '0' after 410 ns,  
		'1' after 424 ns, '0' after 430 ns, 
		'1' after 444 ns, '0' after 450 ns,  
		'1' after 464 ns, '0' after 470 ns, 
		'1' after 484 ns, '0' after 490 ns,
		'1' after 504 ns, '0' after 510 ns,  
		'1' after 524 ns, '0' after 530 ns, 
		'1' after 544 ns, '0' after 550 ns,  
		'1' after 564 ns, '0' after 570 ns, 
		'1' after 584 ns, '0' after 590 ns,
		'1' after 604 ns, '0' after 610 ns,  
		'1' after 624 ns, '0' after 630 ns, 
		'1' after 644 ns, '0' after 650 ns,  
		'1' after 664 ns, '0' after 670 ns, 
		'1' after 684 ns, '0' after 690 ns,
		'1' after 704 ns, '0' after 710 ns,  
		'1' after 724 ns, '0' after 730 ns, 
		'1' after 744 ns, '0' after 750 ns,  
		'1' after 764 ns, '0' after 770 ns, 
		'1' after 784 ns, '0' after 790 ns;
SENSOR_VAGA_SOJA <= '0', 
		'1' after 4 ns, '0' after 10 ns, 
		'1' after 14 ns, '0' after 20 ns, 
		'1' after 24 ns, '0' after 30 ns, 
		'1' after 34 ns, '0' after 40 ns,  
		'1' after 64 ns, '0' after 70 ns, 
		'1' after 74 ns, '0' after 80 ns,
		'1' after 104 ns, '0' after 110 ns, 
		'1' after 114 ns, '0' after 120 ns,  
		'1' after 144 ns, '0' after 150 ns, 
		'1' after 154 ns, '0' after 160 ns, 
		'1' after 184 ns, '0' after 190 ns,
		'1' after 194 ns, '0' after 200 ns,
		'1' after 204 ns, '0' after 210 ns, 
		'1' after 214 ns, '0' after 220 ns, 
		'1' after 224 ns, '0' after 230 ns, 
		'1' after 234 ns, '0' after 240 ns,  
		'1' after 264 ns, '0' after 270 ns, 
		'1' after 274 ns, '0' after 280 ns,
		'1' after 304 ns, '0' after 310 ns, 
		'1' after 314 ns, '0' after 320 ns,  
		'1' after 344 ns, '0' after 350 ns, 
		'1' after 354 ns, '0' after 360 ns, 
		'1' after 384 ns, '0' after 390 ns,
		'1' after 394 ns, '0' after 400 ns,
		'1' after 404 ns, '0' after 410 ns, 
		'1' after 414 ns, '0' after 420 ns, 
		'1' after 424 ns, '0' after 430 ns, 
		'1' after 434 ns, '0' after 440 ns,  
		'1' after 464 ns, '0' after 470 ns, 
		'1' after 474 ns, '0' after 480 ns,
		'1' after 504 ns, '0' after 510 ns, 
		'1' after 514 ns, '0' after 520 ns,  
		'1' after 544 ns, '0' after 550 ns, 
		'1' after 554 ns, '0' after 560 ns, 
		'1' after 584 ns, '0' after 590 ns,
		'1' after 594 ns, '0' after 600 ns,
		'1' after 604 ns, '0' after 610 ns, 
		'1' after 614 ns, '0' after 620 ns, 
		'1' after 644 ns, '0' after 650 ns, 
		'1' after 654 ns, '0' after 660 ns, 
		'1' after 684 ns, '0' after 690 ns,
		'1' after 694 ns, '0' after 700 ns,
		'1' after 704 ns, '0' after 710 ns, 
		'1' after 714 ns, '0' after 720 ns, 
		'1' after 744 ns, '0' after 750 ns, 
		'1' after 754 ns, '0' after 760 ns, 
		'1' after 784 ns, '0' after 790 ns,
		'1' after 794 ns, '0' after 800 ns;
SENSOR_VAGA_ARROZ <= '0', 
		'1' after 4 ns, '0' after 10 ns, 
		'1' after 14 ns, '0' after 20 ns, 
		'1' after 24 ns, '0' after 30 ns, 
		'1' after 34 ns, '0' after 40 ns,  
		'1' after 64 ns, '0' after 70 ns, 
		'1' after 74 ns, '0' after 80 ns,
		'1' after 104 ns, '0' after 110 ns, 
		'1' after 114 ns, '0' after 120 ns,  
		'1' after 144 ns, '0' after 150 ns, 
		'1' after 154 ns, '0' after 160 ns, 
		'1' after 184 ns, '0' after 190 ns,
		'1' after 194 ns, '0' after 200 ns,
		'1' after 204 ns, '0' after 210 ns, 
		'1' after 214 ns, '0' after 220 ns, 
		'1' after 224 ns, '0' after 230 ns, 
		'1' after 234 ns, '0' after 240 ns,  
		'1' after 264 ns, '0' after 270 ns, 
		'1' after 274 ns, '0' after 280 ns,
		'1' after 304 ns, '0' after 310 ns, 
		'1' after 314 ns, '0' after 320 ns,  
		'1' after 344 ns, '0' after 350 ns, 
		'1' after 354 ns, '0' after 360 ns, 
		'1' after 384 ns, '0' after 390 ns,
		'1' after 394 ns, '0' after 400 ns,
		'1' after 404 ns, '0' after 410 ns, 
		'1' after 414 ns, '0' after 420 ns, 
		'1' after 424 ns, '0' after 430 ns, 
		'1' after 434 ns, '0' after 440 ns,  
		'1' after 464 ns, '0' after 470 ns, 
		'1' after 474 ns, '0' after 480 ns,
		'1' after 504 ns, '0' after 510 ns, 
		'1' after 514 ns, '0' after 520 ns,  
		'1' after 544 ns, '0' after 550 ns, 
		'1' after 554 ns, '0' after 560 ns, 
		'1' after 584 ns, '0' after 590 ns,
		'1' after 594 ns, '0' after 600 ns,
		'1' after 604 ns, '0' after 610 ns, 
		'1' after 614 ns, '0' after 620 ns, 
		'1' after 644 ns, '0' after 650 ns, 
		'1' after 654 ns, '0' after 660 ns, 
		'1' after 684 ns, '0' after 690 ns,
		'1' after 694 ns, '0' after 700 ns,
		'1' after 704 ns, '0' after 710 ns, 
		'1' after 714 ns, '0' after 720 ns, 
		'1' after 744 ns, '0' after 750 ns, 
		'1' after 754 ns, '0' after 760 ns, 
		'1' after 784 ns, '0' after 790 ns,
		'1' after 794 ns, '0' after 800 ns;
SENSOR_VAGA_FEIJAO <= '0', 
		'1' after 4 ns, '0' after 10 ns, 
		'1' after 14 ns, '0' after 20 ns, 
		'1' after 24 ns, '0' after 30 ns, 
		'1' after 34 ns, '0' after 40 ns,  
		'1' after 64 ns, '0' after 70 ns, 
		'1' after 74 ns, '0' after 80 ns,
		'1' after 104 ns, '0' after 110 ns, 
		'1' after 114 ns, '0' after 120 ns, 
		'1' after 144 ns, '0' after 150 ns, 
		'1' after 154 ns, '0' after 160 ns, 
		'1' after 184 ns, '0' after 190 ns,
		'1' after 194 ns, '0' after 200 ns,
		'1' after 204 ns, '0' after 210 ns, 
		'1' after 214 ns, '0' after 220 ns, 
		'1' after 224 ns, '0' after 230 ns, 
		'1' after 234 ns, '0' after 240 ns, 
		'1' after 264 ns, '0' after 270 ns, 
		'1' after 274 ns, '0' after 280 ns,
		'1' after 304 ns, '0' after 310 ns, 
		'1' after 314 ns, '0' after 320 ns, 
		'1' after 344 ns, '0' after 350 ns, 
		'1' after 354 ns, '0' after 360 ns, 
		'1' after 384 ns, '0' after 390 ns,
		'1' after 394 ns, '0' after 400 ns,
		'1' after 404 ns, '0' after 410 ns, 
		'1' after 414 ns, '0' after 420 ns, 
		'1' after 424 ns, '0' after 430 ns, 
		'1' after 434 ns, '0' after 440 ns,  
		'1' after 464 ns, '0' after 470 ns, 
		'1' after 474 ns, '0' after 480 ns,
		'1' after 504 ns, '0' after 510 ns, 
		'1' after 514 ns, '0' after 520 ns, 
		'1' after 544 ns, '0' after 550 ns, 
		'1' after 554 ns, '0' after 560 ns, 
		'1' after 584 ns, '0' after 590 ns,
		'1' after 594 ns, '0' after 600 ns,
		'1' after 604 ns, '0' after 610 ns, 
		'1' after 614 ns, '0' after 620 ns, 
		'1' after 644 ns, '0' after 650 ns, 
		'1' after 654 ns, '0' after 660 ns, 
		'1' after 684 ns, '0' after 690 ns,
		'1' after 694 ns, '0' after 700 ns,
		'1' after 704 ns, '0' after 710 ns, 
		'1' after 714 ns, '0' after 720 ns, 
		'1' after 744 ns, '0' after 750 ns, 
		'1' after 754 ns, '0' after 760 ns, 
		'1' after 784 ns, '0' after 790 ns,
		'1' after 794 ns, '0' after 800 ns;
		
PESO_BRUTO <= "00000000000010011100010000000",
					"00000000000011000011010100000" after 275 ns,
					"00000000000010001000101110000" after 515 ns;
PESO_CAMINHAO <= "00000000000000010011100010000",
						"00000000000001010010000010000" after 275 ns,
						"00000000000000110100101111000" after 515 ns;
TIPO_GRAO <= "10",
					"01" after 275 ns,
					"11" after 515 ns;		
--PESO_BRUTO <= std_logic_vector(to_unsigned(80000, 32)),
--					std_logic_vector(to_unsigned(100000, 32)) after 200 ns,
--					std_logic_vector(to_unsigned(70000, 32)) after 400 ns;
--PESO_CAMINHAO <= std_logic_vector(to_unsigned(10000, 32)),
--						std_logic_vector(to_unsigned(42000, 32)) after 200 ns,
--						std_logic_vector(to_unsigned(27000, 32)) after 400 ns;
--TIPO_GRAO <= std_logic_vector(to_unsigned(2, 2)),
--					std_logic_vector(to_unsigned(1, 2)) after 200 ns,
--					std_logic_vector(to_unsigned(3, 2)) after 400 ns;
end teste;